module alu_controller (
    ia, ib, func,
    oa
);

input   [7:0] ia;
input   [7:0] ib;
input   [3:0] func;
output reg [7:0] oa;

alu_8bit U0_alu_8bit(

)
    
endmodule